dncdsn

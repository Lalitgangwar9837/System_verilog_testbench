https://www.edaplayground.com/x/JnjQ

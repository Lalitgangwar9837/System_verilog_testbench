
interface bus ;
  logic [3:0] sum,a,b;
  logic carry;
  
  
endinterface
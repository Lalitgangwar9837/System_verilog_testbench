interface intf;
  logic a;
  logic b;
  logic carry_in;
  logic sum;
  logic carry;
  
endinterface
interface intf(input logic clk, rst);
  logic [3:0]cnt;
endinterface
